module comparador(
   input logic [6:0] data_paridad, 
   output logic [6:0] comparacion);
endmodule