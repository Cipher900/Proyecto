`timescale 1ns/1ns

module module_top_tb;
endmodule